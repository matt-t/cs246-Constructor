0
6 5 4 2 5 r 32 0 h 1 B 21 H
0 1 2 2 3 r h 3 T 19 T 37 T
10 10 10 10 10 r h 5 B 11 B 24 T 
3 2 1 0 1 r h 50 B 36 B
2 4 5 7 4 6 1 8 1 8 3 5 2 5 0 11 3 2 4 3 4 4 3 9 0 10 4 11 2 10 0 3 2 6 3 9 4 5 