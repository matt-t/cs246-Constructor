2
10 10 10 10 10 r h 5 B 21 H 24 T 33 B
3 2 1 0 1 r h 50 B 36 B
2 10 10 10 0 r h 3 T 26 T 37 T
3 2 5 1 7 r 0 h 1 B 11 H 34 B
5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 5 7 