45
2 2 1 0 5 r 1 3 6 14 22 31 h 2 B 0 B
0 0 0 2 2 r 7 10 h 4 B 27 B
0 2 0 5 20 r h 13 B 25 B
0 2 0 5 0 r h 15 B 17 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
