0
6 5 4 2 5 r 32 0 h 1 B 21 H
0 1 2 2 3 r h 3 T 19 T 37 T
10 10 10 10 10 r h 5 B 11 B 24 T 
3 2 1 0 1 r h 
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
