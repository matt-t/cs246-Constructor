0
0 0 0 0 0 r h 1 B 20 B
0 0 0 1 0 r h 3 B 30 B
0 0 0 0 0 r h 5 B 50 B
0 0 0 0 0 r h 7 B 9 B
2 4 5 7 4 6 1 8 1 8 3 5 2 5 0 11 3 2 4 3 4 4 3 9 0 10 4 11 2 10 0 3 2 6 3 9 4 5
