3
1 2 3 4 5 r 2 7 h 1 B 11 B 36 H
0 1 2 2 3 r h 3 B 26 H 37 T
10 9 8 7 6 r h 5 B 21 H 24 T 33 B
0 0 0 0 11 r h 50 B 34 B
2 4 5 7 4 6 1 8 1 8 3 5 2 5 0 11 3 2 4 3 4 4 3 9 0 10 4 11 2 10 0 3 2 6 3 9 4 5 
11
