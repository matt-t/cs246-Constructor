1
10 11 10 9 9 r 3 h 2 B 29 H
10 10 10 10 10 r h 4 T 27 B
10 11 10 10 10 r h 13 B 25 B
10 10 10 11 10 r h 15 B 17 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
1
