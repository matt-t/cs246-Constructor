0
3 3 3 5 3 r 38 47 43 h 25 T 30 B 37 T
0 0 0 0 0 r 56 48 64 h 32 H 44 B
11 0 0 0 0 r 24 50 33 41 h 16 H 40 B
0 0 3 0 0 r 27 32 h 20 H 27 H
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
3
