<<<<<<< HEAD
0
0 0 0 0 0 r h 1 B 20 B
0 0 0 1 0 r h 3 B 30 B
0 0 0 0 0 r h 5 B 50 B
0 0 0 0 0 r h 7 B 9 B
2 4 5 7 4 6 1 8 1 8 3 5 2 5 0 11 3 2 4 3 4 4 3 9 0 10 4 11 2 10 0 3 2 6 3 9 4 5
=======
4
0 1 2 2 3 r 2 7 h 1 B 11 B 36 H
0 1 1 0 4 r h 3 B 26 H 37 T
4 6 4 2 7 r h 5 B 21 H 24 T 33 B
1 0 0 0 6 r h 34 B 50 B
2 4 5 7 4 6 1 8 1 8 3 5 2 5 0 11 3 2 4 3 4 4 3 9 0 10 4 11 2 10 0 3 2 6 3 9 4 5
9
>>>>>>> 299172aded00b7c532955311275e3998be9c61c2
