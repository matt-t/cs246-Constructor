10
1 0 0 0 0 r h 2 B 29 B
2 0 0 0 3 r h 4 B 27 B
0 2 0 1 0 r h 13 B 25 B
1 0 0 0 0 r h 15 B 17 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
