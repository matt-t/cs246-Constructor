1
10 10 10 10 10 r h
9 9 9 9 8 r 71 70 h 53 B
10 10 10 10 10 r h
10 10 10 10 10 r h
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
0